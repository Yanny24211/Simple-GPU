LIBRARY ieee; 
USE ieee.std_logic_1164.all;

ENTITY modsseg IS 
	PORT ( 
			bcd 	: 	IN STD_LOGIC_VECTOR(3 DOWNTO 0) ; 
			yn	: 	OUT STD_LOGIC_VECTOR(0 TO 6)
			);
END modsseg;

ARCHITECTURE Behavior OF modsseg IS 
BEGIN 
	PROCESS ( bcd ) 
	BEGIN
		CASE bcd IS
			
			WHEN "0000"  => yn <= "0111011"; 
			WHEN "0001"	 => yn <= "0010101";
			WHEN OTHERS  => yn <= "-------";
		END CASE; 
	END PROCESS;
END Behavior ;